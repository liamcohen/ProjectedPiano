`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Zoe Klawans
// 
// Create Date:    15:24:29 11/28/2017 
// Design Name: 
// Module Name:    keystoning 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module keystoning(
    input clk,
    input reset,
	 input [10:0] hcount,
	 input [9:0] vcount,
	 input hsync,
	 input vsync,
	 input blank,
	 input [16:0] key_num,
	 input note_ready,
	 input [1:0] state,
	 
	 output phsync,
	 output pvsync,
	 output pblank,
    output [23:0] keystoned_pixel
    );
	
	parameter WHITE_KEY_WIDTH = 99;
	parameter SPACE = 4;
	parameter PIANO_MIDDLE = (5 * WHITE_KEY_WIDTH) + (4 * SPACE) + 2;
	parameter BOARD_HEIGHT = 10'd768;
	parameter KEY_START_VERTICAL = BOARD_HEIGHT >> 2;
   parameter WHITE_KEY_HEIGHT = BOARD_HEIGHT >> 2;
	parameter PIANO_LENGTH = (10 * WHITE_KEY_WIDTH) + (9 * SPACE);
	parameter PIANO_HALF = PIANO_LENGTH >> 1;
	parameter BLACK = 24'h00_00_00;
	parameter RED = 24'hFF_00_00;
	parameter GREEN = 24'h00_FF_00;
	
	reg [10:0] phcount;
	reg [9:0] pvcount;
	reg signed [10:0] x;
	wire [23:0] temp_pixel;
	
	always @(posedge clk)
	begin
		
		x <= hcount - PIANO_MIDDLE;
//		if (x < 0) phcount <= hcount - (((vcount - KEY_START_VERTICAL) * (x * -1)) >> 9);
//		else phcount <= hcount - (((vcount - KEY_START_VERTICAL) * (x * -1)) >> 9);
		phcount <= hcount - (((vcount - KEY_START_VERTICAL) * (x * -1)) >> 10);
		
	end
	
	piano p(.vclock(clk), .reset(reset), .hcount(phcount), .vcount(vcount),
			.hsync(hsync), .vsync(vsync), .blank(blank), .key_num(key_num),
			.note_ready(note_ready), .state(state), .phsync(phsync), .pvsync(pvsync),
			.pblank(pblank), .pixel(temp_pixel));
	
	assign keystoned_pixel = (hcount < 2) ? BLACK : temp_pixel;
		
endmodule
